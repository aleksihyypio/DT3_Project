
package apb_env_pkg;

`ifndef SYNTHESIS
   
`include "uvm_macros.svh"

   import uvm_pkg::*;
   import apb_pkg::*;
   import audioport_pkg::*;
   
`include "apb_transaction.svh"
`include "apb_driver.svh"
`include "apb_monitor.svh"
`include "apb_analyzer.svh"
`include "apb_sequencer.svh"
`include "apb_agent_config.svh"   
`include "apb_agent.svh"
`include "apb_env.svh"

`endif //  `ifndef SYNTHESIS
   
endpackage

   


