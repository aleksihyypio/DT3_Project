//
//  audioport.sv: Top-level module of audioport design.
//

`include "audioport.svh"

import audioport_pkg::*;

module audioport
  
  (input logic clk,
   input logic 	       rst_n,
   input logic 	       mclk,
   // APB interface
   input logic 	       PSEL,
   input logic 	       PENABLE,
   input logic 	       PWRITE,
   input logic [31:0]  PADDR,
   input logic [31:0]  PWDATA,
   output logic [31:0] PRDATA,
   output logic        PREADY,
   output logic        PSLVERR,
   // Interrupt request
   output logic        irq_out,
   // Audio outputs
   output logic        ws_out,
   output logic        sck_out, 
   output logic        sdo_out,
   // Test signals
   input logic 	       test_mode_in,
   input logic 	       scan_en_in
   );

   /////////////////////////////////////////////////////////////////////////////
   // Internal variables
   /////////////////////////////////////////////////////////////////////////////
   

   
   /////////////////////////////////////////////////////////////////////////////
   // control_unit instantiation
   /////////////////////////////////////////////////////////////////////////////
   

   /////////////////////////////////////////////////////////////////////////////
   // dsp_unit instantiation
   /////////////////////////////////////////////////////////////////////////////
   

   /////////////////////////////////////////////////////////////////////////////
   // cdc_unit instantiation
   /////////////////////////////////////////////////////////////////////////////
   

   /////////////////////////////////////////////////////////////////////////////
   // i2s_unit instantiation
   /////////////////////////////////////////////////////////////////////////////
   

endmodule


